library verilog;
use verilog.vl_types.all;
entity bcd_add_test is
end bcd_add_test;
