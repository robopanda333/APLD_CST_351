library verilog;
use verilog.vl_types.all;
entity test_ClkDiv is
end test_ClkDiv;
