library verilog;
use verilog.vl_types.all;
entity test_alu_top_level is
end test_alu_top_level;
